library IEEE;
use IEEE.STD_LOGIC_1164.all;

package constants is

constant CLOCK_DIVIDER_1MS: integer:= 106250;
 

end constants;
